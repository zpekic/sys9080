----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 09/24/2017 10:11:13 AM
-- Design Name: 
-- Module Name: Am25LS377 - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: https://datasheet.datasheetarchive.com/originals/scans/Scans-001/Scans-0034821.pdf
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Am25LS377 is
    Port ( clk : in STD_LOGIC;
           nE : in STD_LOGIC;
           d : in STD_LOGIC_VECTOR (7 downto 0);
           q : out STD_LOGIC_VECTOR (7 downto 0));
end Am25LS377;

architecture Behavioral of Am25LS377 is

begin

update_q: process(clk, nE, d)
begin
	if (nE = '0') then
		if (rising_edge(clk)) then
        q <= d;
		end if;
	end if;
end process;

end Behavioral;
